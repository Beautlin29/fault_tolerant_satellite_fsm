module top(I1, I2, I3, C1, C2, Sel, N1, N2);
    input [86:1]Sel;
    input I1, I2, I3, C1, C2;
    output N1, N2;
    wire [14:1]x;
    wire [10:1]y;
    wire [5:1]z;
    wire [4:1]zz;

    //Sel = 86'b0101_0110_0010_011_0101_0001_0111_0100_100_1_0101_0110_1000_011_0001_0010_0011_011_0101_0010_0011_1001_100_1;


    //PE1 --> ~I1.~I2.I3
    mux_16_1 a1 (x[1], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[86:83]);
    mux_16_1 a2 (x[2], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[82:79]);
    mux_16_1 a3 (x[3], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[78:75]);

    and_3 b1 (x[1], x[2], x[3], y[1]);
    or_3 c1 (x[1], x[2], x[3], y[2]);

    mux_8_1 aa1 (z[1], x[1], x[2], x[3], y[1], y[2], 1'bx, 1'bx, 1'bx, Sel[74:72]);


    //PE2 --> ~I1.I2.~I3.C2
    mux_16_1 a4 (x[4], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[71:68]);
    mux_16_1 a5 (x[5], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[67:64]);
    mux_16_1 a6 (x[6], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[63:60]);
    mux_16_1 a7 (x[7], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[59:56]);

    and_4 b2 (x[4], x[5], x[6], x[7], y[3]);
    or_4 c2 (x[4], x[5], x[6], x[7], y[4]);

    mux_8_1 aa2 (z[2], x[4], x[5], x[6], x[7], y[3], y[4], 1'bx, 1'bx, Sel[55:53]);

    //N1
    and_2 b3 (z[1], z[2], zz[1]);
    or_2 c3 (z[1], z[2], zz[2]);
    mux_2_1 aaa1 (N1, zz[1], zz[2], Sel[52]);

    //--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------//

    //PE3 --> ~I1.~I2.~C1
    mux_16_1 a8 (x[8], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[51:48]);
    mux_16_1 a9 (x[9], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[47:44]);
    mux_16_1 a10 (x[10], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[43:40]);

    and_3 b4 (x[8], x[9], x[10], y[5]);
    or_3 c4 (x[8], x[9], x[10], y[6]);

    mux_8_1 aa3 (z[3], x[8], x[9], x[10], y[5], y[6], 1'bx, 1'bx, 1'bx, Sel[39:37]);


    //PE4 --> C1.I2.I3
    mux_16_1 a11 (x[11], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[36:33]);
    mux_16_1 a12 (x[12], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[32:29]);
    mux_16_1 a13 (x[13], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[28:23]);

    and_3 b5 (x[11], x[12], x[13], y[7]);
    or_3 c5 (x[11], x[12], x[13], y[8]);

    mux_8_1 aa4 (z[4], x[11], x[12], x[13], y[7], y[8], 1'bx, 1'bx, 1'bx,  Sel[24:21]);


    //PE5 --> ~I1.I3.C1.~C2
    mux_16_1 a14 (x[14], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[20:17]);
    mux_16_1 a15 (x[15], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[16:13]);
    mux_16_1 a16 (x[16], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[12:9]);
    mux_16_1 a17 (x[17], I1, I2, I3, C1, C2, ~I1, ~I2, ~I3, ~C1, ~C2, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, 1'bx, Sel[8:5]);

    and_4 b6 (x[14], x[15], x[16], x[17], y[9]);
    or_4 c6 (x[14], x[15], x[16], x[17], y[10]);

    mux_8_1 aa5 (z[5], x[14], x[15], x[16], x[17], y[9], y[10], 1'bx, 1'bx, Sel[4:2]);

    //N2
    and_3 b7 (z[3], z[4], z[5], zz[3]);
    or_3 c7 (z[3], z[4], z[5], zz[4]);
    mux_2_1 aaa2 (N2, zz[3], zz[4], Sel[1]);


endmodule
